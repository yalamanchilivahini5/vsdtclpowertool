* source INV
M_M1         OUT N14434 0 0 NMOS  
+ L=.18u  
+ W=.76u         
M_M2         OUT N14434 net net PMOS  
+ L=.18u  
+ W=1.8u         
V_V1         VDD 0 1.8Vdc
V_V2         N14434 0  
+PULSE 1.8V 0V 0ns 1ns 1ns 2us 4us
C_C1         0 OUT  20p   
Vnet         VDD net 0Vdc
 
Fnet 0 netl Vnet 1.0
Cnet netl 0 1.111u
Rnet netl 0 111100.0k 
 
.MODEL PMOS PMOS
.MODEL NMOS NMOS  

.tran 2e-0 20e-6 2e-6 uic
.control
run
plot V(netl)
wrdata outinverter.txt V(netl)
.endc
.end